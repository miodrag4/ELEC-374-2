module Memory_Subsystem();

endmodule
