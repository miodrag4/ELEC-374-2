module Decoder4to16(     
input [3:0] Din,    
output reg [15:0] Dout 
);

always @(*) begin   
	case (Din)
		4'b0000: Dout = 16'b0000000000000001;         
		4'b0001: Dout = 16'b0000000000000010;         
		4'b0010: Dout = 16'b0000000000000100;         
		4'b0011: Dout = 16'b0000000000001000;         
		4'b0100: Dout = 16'b0000000000010000;         
		4'b0101: Dout = 16'b0000000000100000;         
		4'b0110: Dout = 16'b0000000001000000;         
		4'b0111: Dout = 16'b0000000010000000;         
		4'b1000: Dout = 16'b0000000100000000;         
		4'b1001: Dout = 16'b0000001000000000;         
		4'b1010: Dout = 16'b0000010000000000;         
		4'b1011: Dout = 16'b0000100000000000;         
		4'b1100: Dout = 16'b0001000000000000;         
		4'b1101: Dout = 16'b0010000000000000;         
		4'b1110: Dout = 16'b0100000000000000;         
		4'b1111: Dout = 16'b1000000000000000;
		default Dout = 16'bx;
		endcase 
end 
endmodule
